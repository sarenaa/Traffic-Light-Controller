package light_package;

typedef enum logic[1:0] {red,yellow,green} colors;

endpackage